/****************************************************************

Copyright (c) 2018- Stanford University. All rights reserved.

The information and source code contained herein is the 
property of Stanford University, and may not be disclosed or
reproduced in whole or in part without explicit written 
authorization from Stanford University. Contact bclim@stanford.edu for details.

* Filename   : buck_core.v
* Author     : Byongchan Lim (bclim@stanford.edu)
* Description: Output driver of a buck converter

* Note       :

* Revision   :
  - 7/26/2016: First release

****************************************************************/


module buck_core #(
  parameter rp = 0.4,
  parameter CL = 1e-12, 
  parameter L = 1e-09, 
  parameter RL = 100, 
  parameter etol = 0.001 // error tolerance of PWL approximation
) (
  input din, // up & dn driver's input
  `input_pwl vddh, vgnd,     // power & ground
  `output_real swout,  // switch output signal for feedback
  `output_pwl so
);

`get_timeunit
PWLMethod pm=new;

real si;
real poler, polei;
real p1, p2;
real prelax;
real sqterm;
reg sqterm_isreal=1'b0;
reg up_or_dn=1'b1;  // din_up | din_dn 
reg up_or_dn_prev=1'b0;

always @(si) swout = si;

// pole location
initial begin
  sqterm = CL**2*RL**2*rp**2 - 4*CL*L*RL**2 - 2*CL*L*RL*rp + L**2;
  if (sqterm >=0) begin
    p2 = 0.5*(CL*RL*rp + L)/(CL*L*RL) - 0.5*sqrt(sqterm)/(CL*L*RL); 
    p1 = 0.5*(CL*RL*rp + L)/(CL*L*RL) + 0.5*sqrt(sqterm)/(CL*L*RL); 
    sqterm_isreal = 1'b1;
  end
  else begin
    poler = 0.5*(CL*RL*rp + L)/(CL*L*RL);
    polei = 0.5*sqrt(-1*(CL**2*RL**2*rp**2 - 4*CL*L*RL**2 - 2*CL*L*RL*rp + L**2))/(CL*L*RL);
    sqterm_isreal = 1'b0;
  end
end

always @(din or `pwl_event(vddh) or `pwl_event(vgnd)) begin
  // assertion
  if (~din) si = pm.eval(vddh, `get_time);
  else si = pm.eval(vgnd, `get_time);
end


/***************************************************************
 Generated by PWL analog filter model generator in SystemVerilog

 Copyright (c) 2014- by Byong Chan Lim. All rights reserved.

 The information and source code contained herein is the property
 of Byong Chan Lim, and may not be disclosed or reproduced
 in whole or in part without explicit written authorization from
 Byong Chan Lim.
 ***************************************************************/


// wires
event wakeup;  // event signal
real t0;  // time offset
real t_cur;   // current time
real dTr;  // time interval of PWL waveform
time dT=1;
time dTm, t_prev;
reg event_in=1'b0;

real si_at_t0;  // 
real so_cur; // current output signal value
real so_prev; // previous output signal value
real so_nxt;  // so at (t_cur+dT) for pwl output data
real yo0;  // output signal value offset (so_cur at t0)
real yo1;  // first derivative y'(0)
real xi0;  // initial state of input
real xi1;  // initial state of first derivative of input

real so_slope; // so slope

initial so = '{0,0,0};

reg dum;

always @(si) begin
  t0 = `get_time;
  so_cur = pm.eval(so, t0);
  si_at_t0 = si;
  yo0 = so_cur;
  yo1 = so.b;
  xi0 = si;

  t_prev = $realtime;
  dT = 0;
  ->> wakeup;
end

always @(wakeup) begin
  dTm = $realtime - t_prev;
  
  if (dT==dTm) begin
    t_prev = $realtime;
    t_cur = `get_time;
    so_cur = pm.eval(so, t_cur);
    
    // calculate next time step (dTr)
    dTr = calculate_Tintv_buck(etol, t_cur-t0, si_at_t0, xi0, xi1, yo0, yo1  );
    //dTr = min(1,max(TU,dTr));
    dT = time'(dTr/TU);

    so_nxt = fn_buck(t_cur-t0+dTr, si_at_t0, xi0, xi1, yo0, yo1  );
    so_slope = (so_nxt-so_cur)/dTr;
    so = pm.write(so_cur, so_slope, t_cur);

    // schedule next event
    if (so_slope != 0) ->> #(dT) wakeup;
  end

end

/*******************************************
  Response function, its 1st/2nd derivatives
*******************************************/

function real fn_buck;
input real t; 
input real si; 
input real xi0, xi1, yo0, yo1  ;
begin
  if (up_or_dn) begin
    if (sqterm_isreal)
      return si/(CL*L*p1*p2) + ((CL*L*p1*p2*yo0 + CL*L*p2*yo1 - si)/(CL*L*p2*(p1 - p2)))*exp(-1.0*t/(1/p2)) + (-(CL*L*p1*p2*yo0 + CL*L*p1*yo1 - si)/(CL*L*p1*(p1 - p2)))*exp(-1.0*t/(1/p1));
    else
      return si/(CL*L*polei**2 + CL*L*poler**2) - (-CL*L*polei**2*yo0*cos(polei*t) - CL*L*polei*yo1*sin(polei*t) - CL*L*poler**2*yo0*cos(polei*t) - CL*L*poler*yo1*cos(polei*t) + si*cos(polei*t))*exp(-poler*t)/(2*CL*L*(polei**2 + poler**2)) + (CL*L*polei**2*yo0*cos(polei*t) + CL*L*polei*yo1*sin(polei*t) + CL*L*poler**2*yo0*cos(polei*t) + CL*L*poler*yo1*cos(polei*t) - si*cos(polei*t))*exp(-poler*t)/(2*CL*L*(polei**2 + poler**2)) + poler*(CL*L*polei**2*yo0*sin(polei*t) - CL*L*polei*yo1*cos(polei*t) + CL*L*poler**2*yo0*sin(polei*t) + CL*L*poler*yo1*sin(polei*t) - si*sin(polei*t))*exp(-poler*t)/(CL*L*polei*(polei**2 + poler**2));
  end
  else
    return yo0*exp(-prelax*t);
end
endfunction

function real f2max_buck;
input real t; 
input real si; 
input real xi0, xi1, yo0, yo1  ;
begin
  if (up_or_dn) begin
    if (sqterm_isreal)
      return abs((CL*L*p1*p2*yo0 + CL*L*p2*yo1 - si)/(CL*L*p2*(p1 - p2)))*p2**2*exp(-p2*t) + abs(-(CL*L*p1*p2*yo0 + CL*L*p1*yo1 - si)/(CL*L*p1*(p1 - p2)))*p1**2*exp(-p1*t);
    else 
      return abs((-polei**2*(CL*L*polei**2*yo0*cos(polei*t) + CL*L*polei*yo1*sin(polei*t) + CL*L*poler**2*yo0*cos(polei*t) + CL*L*poler*yo1*cos(polei*t) - si*cos(polei*t)) + polei*poler*(CL*L*polei**2*yo0*sin(polei*t) - CL*L*polei*yo1*cos(polei*t) + CL*L*poler**2*yo0*sin(polei*t) + CL*L*poler*yo1*sin(polei*t) - si*sin(polei*t)) - poler**2*(CL*L*polei**2*yo0*cos(polei*t) + CL*L*polei*yo1*sin(polei*t) + CL*L*poler**2*yo0*cos(polei*t) + CL*L*poler*yo1*cos(polei*t) - si*cos(polei*t)) + poler**3*(CL*L*polei**2*yo0*sin(polei*t) - CL*L*polei*yo1*cos(polei*t) + CL*L*poler**2*yo0*sin(polei*t) + CL*L*poler*yo1*sin(polei*t) - si*sin(polei*t))/polei)*exp(-poler*t)/(CL*L*(polei**2 + poler**2)));
  end
  else
    return abs(yo0)*prelax**2*exp(-prelax*t);
end
endfunction

/*************************************
  Caluating Tintv
*************************************/

function real calculate_Tintv_buck;
input real etol, t; 
input real si; 
input real xi0, xi1, yo0, yo1  ;
real abs_f2max;
real calcT;
begin
  abs_f2max = f2max_buck(t, si, xi0, xi1, yo0, yo1  );
  calcT = sqrt(8.0*etol/abs_f2max);
  return max(TU,min(1.0,calcT));
  //return sqrt(8.0*etol/abs_f2max); 
end
endfunction

endmodule
