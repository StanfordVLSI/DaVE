../../../include/pwlgen.vh