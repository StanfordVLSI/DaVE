// dummy module

module comparator (
  input real vinp, vinn,
  output real voutp, voutn,
  input pdn, clk_preamp, clk_latch,
  output out, outb
);

endmodule
